module ctrl (clk, reset);

  

endmodule